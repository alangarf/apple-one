module ukprom(clk, adr, data);
	input clk;
	input [9:0] adr;
	output [3:0] data;
	reg [3:0] data;
	always @(posedge clk) begin
		case (adr)
			10'h000: data <= 4'h1;
			10'h001: data <= 4'h9;
			10'h002: data <= 4'h0;
			10'h003: data <= 4'h0;
			10'h004: data <= 4'he;
			10'h005: data <= 4'h9;
			10'h006: data <= 4'h2;
			10'h007: data <= 4'h8;
			10'h008: data <= 4'h8;
			10'h009: data <= 4'h0;
			10'h00a: data <= 4'h0;
			10'h00b: data <= 4'h1;
`ifdef SIM
			10'h00c: data <= 4'h2;
			10'h00d: data <= 4'h0;
`else
			10'h00c: data <= 4'h8;
			10'h00d: data <= 4'hc;
`endif
			10'h00e: data <= 4'h0;
			10'h00f: data <= 4'h0;
			10'h010: data <= 4'he;
			10'h011: data <= 4'hb;
			10'h012: data <= 4'h4;
			10'h013: data <= 4'h0;
			10'h014: data <= 4'h4;
			10'h015: data <= 4'h1;
`ifdef SIM
			10'h016: data <= 4'h1;
			10'h017: data <= 4'h0;
`else
			10'h016: data <= 4'ha;
			10'h017: data <= 4'h0;
`endif
			10'h018: data <= 4'he;
			10'h019: data <= 4'hb;
			10'h01a: data <= 4'h6;
			10'h01b: data <= 4'h0;
			10'h01c: data <= 4'h7;
			10'h01d: data <= 4'h1;
`ifdef SIM
			10'h01e: data <= 4'h1;
			10'h01f: data <= 4'h0;
`else
			10'h01e: data <= 4'h8;
			10'h01f: data <= 4'h2;
`endif
			10'h020: data <= 4'he;
			10'h021: data <= 4'h4;
			10'h022: data <= 4'h4;
			10'h023: data <= 4'h6;
			10'h024: data <= 4'h6;
			10'h025: data <= 4'h7;
			10'h026: data <= 4'hb;
			10'h027: data <= 4'h8;
			10'h028: data <= 4'h0;
			10'h029: data <= 4'he;
			10'h02a: data <= 4'h5;
			10'h02b: data <= 4'h6;
			10'h02c: data <= 4'h5;
			10'h02d: data <= 4'h6;
			10'h02e: data <= 4'h5;
			10'h02f: data <= 4'h6;
			10'h030: data <= 4'h5;
			10'h031: data <= 4'h5;
			10'h032: data <= 4'h5;
			10'h033: data <= 4'h6;
			10'h034: data <= 4'h6;
			10'h035: data <= 4'h6;
			10'h036: data <= 4'h5;
			10'h037: data <= 4'h5;
			10'h038: data <= 4'h6;
			10'h039: data <= 4'h5;
			10'h03a: data <= 4'h6;
			10'h03b: data <= 4'h5;
			10'h03c: data <= 4'h6;
			10'h03d: data <= 4'h5;
			10'h03e: data <= 4'h6;
			10'h03f: data <= 4'h5;
			10'h040: data <= 4'h6;
			10'h041: data <= 4'h5;
			10'h042: data <= 4'h6;
			10'h043: data <= 4'h5;
			10'h044: data <= 4'h6;
			10'h045: data <= 4'h5;
			10'h046: data <= 4'h5;
			10'h047: data <= 4'h6;
			10'h048: data <= 4'h5;
			10'h049: data <= 4'h6;
			10'h04a: data <= 4'h4;
			10'h04b: data <= 4'h4;
			10'h04c: data <= 4'h6;
			10'h04d: data <= 4'h6;
			10'h04e: data <= 4'h5;
			10'h04f: data <= 4'h6;
			10'h050: data <= 4'h5;
			10'h051: data <= 4'h6;
			10'h052: data <= 4'h5;
			10'h053: data <= 4'h6;
			10'h054: data <= 4'h5;
			10'h055: data <= 4'h5;
			10'h056: data <= 4'h5;
			10'h057: data <= 4'h5;
			10'h058: data <= 4'h6;
			10'h059: data <= 4'h5;
			10'h05a: data <= 4'h6;
			10'h05b: data <= 4'h5;
			10'h05c: data <= 4'h5;
			10'h05d: data <= 4'h5;
			10'h05e: data <= 4'h6;
			10'h05f: data <= 4'h5;
			10'h060: data <= 4'h6;
			10'h061: data <= 4'h5;
			10'h062: data <= 4'h6;
			10'h063: data <= 4'h5;
			10'h064: data <= 4'h6;
			10'h065: data <= 4'h5;
			10'h066: data <= 4'h5;
			10'h067: data <= 4'h6;
			10'h068: data <= 4'h6;
			10'h069: data <= 4'h5;
			10'h06a: data <= 4'h6;
			10'h06b: data <= 4'h5;
			10'h06c: data <= 4'h6;
			10'h06d: data <= 4'h5;
			10'h06e: data <= 4'h5;
			10'h06f: data <= 4'h6;
			10'h070: data <= 4'h5;
			10'h071: data <= 4'h6;
			10'h072: data <= 4'h5;
			10'h073: data <= 4'h6;
			10'h074: data <= 4'h5;
			10'h075: data <= 4'h6;
			10'h076: data <= 4'h5;
			10'h077: data <= 4'h6;
			10'h078: data <= 4'h5;
			10'h079: data <= 4'h6;
			10'h07a: data <= 4'h5;
			10'h07b: data <= 4'h6;
			10'h07c: data <= 4'h5;
			10'h07d: data <= 4'h6;
			10'h07e: data <= 4'h5;
			10'h07f: data <= 4'h6;
			10'h080: data <= 4'h5;
			10'h081: data <= 4'h6;
			10'h082: data <= 4'h5;
			10'h083: data <= 4'h6;
			10'h084: data <= 4'h5;
			10'h085: data <= 4'h6;
			10'h086: data <= 4'h5;
			10'h087: data <= 4'h6;
			10'h088: data <= 4'h5;
			10'h089: data <= 4'h6;
			10'h08a: data <= 4'h5;
			10'h08b: data <= 4'h6;
			10'h08c: data <= 4'h5;
			10'h08d: data <= 4'h6;
			10'h08e: data <= 4'h5;
			10'h08f: data <= 4'h6;
			10'h090: data <= 4'h5;
			10'h091: data <= 4'h6;
			10'h092: data <= 4'h5;
			10'h093: data <= 4'h6;
			10'h094: data <= 4'h5;
			10'h095: data <= 4'h6;
			10'h096: data <= 4'h5;
			10'h097: data <= 4'h6;
			10'h098: data <= 4'h5;
			10'h099: data <= 4'h6;
			10'h09a: data <= 4'h5;
			10'h09b: data <= 4'h6;
			10'h09c: data <= 4'h5;
			10'h09d: data <= 4'h6;
			10'h09e: data <= 4'h6;
			10'h09f: data <= 4'h6;
			10'h0a0: data <= 4'h5;
			10'h0a1: data <= 4'h5;
			10'h0a2: data <= 4'h6;
			10'h0a3: data <= 4'h6;
			10'h0a4: data <= 4'h6;
			10'h0a5: data <= 4'h6;
			10'h0a6: data <= 4'h6;
			10'h0a7: data <= 4'h5;
			10'h0a8: data <= 4'h5;
			10'h0a9: data <= 4'h6;
			10'h0aa: data <= 4'h5;
			10'h0ab: data <= 4'h5;
			10'h0ac: data <= 4'h6;
			10'h0ad: data <= 4'h5;
			10'h0ae: data <= 4'h4;
			10'h0af: data <= 4'h4;
			10'h0b0: data <= 4'h6;
			10'h0b1: data <= 4'h6;
			10'h0b2: data <= 4'h7;
			10'h0b3: data <= 4'h1;
			10'h0b4: data <= 4'h0;
			10'h0b5: data <= 4'h4;
			10'h0b6: data <= 4'h2;
			10'h0b7: data <= 4'hd;
			10'h0b8: data <= 4'h1;
			10'h0b9: data <= 4'h8;
			10'h0ba: data <= 4'h0;
			10'h0bb: data <= 4'h0;
			10'h0bc: data <= 4'h8;
			10'h0bd: data <= 4'he;
			10'h0be: data <= 4'h2;
			10'h0bf: data <= 4'hb;
			10'h0c0: data <= 4'hf;
			10'h0c1: data <= 4'h2;
			10'h0c2: data <= 4'h0;
			10'h0c3: data <= 4'h0;
			10'h0c4: data <= 4'h5;
			10'h0c5: data <= 4'h6;
			10'h0c6: data <= 4'h5;
			10'h0c7: data <= 4'h6;
			10'h0c8: data <= 4'h5;
			10'h0c9: data <= 4'h6;
			10'h0ca: data <= 4'h5;
			10'h0cb: data <= 4'h5;
			10'h0cc: data <= 4'h5;
			10'h0cd: data <= 4'h6;
			10'h0ce: data <= 4'h5;
			10'h0cf: data <= 4'h5;
			10'h0d0: data <= 4'h6;
			10'h0d1: data <= 4'h6;
			10'h0d2: data <= 4'h6;
			10'h0d3: data <= 4'h5;
			10'h0d4: data <= 4'h6;
			10'h0d5: data <= 4'h5;
			10'h0d6: data <= 4'h6;
			10'h0d7: data <= 4'h5;
			10'h0d8: data <= 4'h6;
			10'h0d9: data <= 4'h5;
			10'h0da: data <= 4'h6;
			10'h0db: data <= 4'h5;
			10'h0dc: data <= 4'h6;
			10'h0dd: data <= 4'h5;
			10'h0de: data <= 4'h6;
			10'h0df: data <= 4'h5;
			10'h0e0: data <= 4'h5;
			10'h0e1: data <= 4'h6;
			10'h0e2: data <= 4'h5;
			10'h0e3: data <= 4'h6;
			10'h0e4: data <= 4'h4;
			10'h0e5: data <= 4'h4;
			10'h0e6: data <= 4'h6;
			10'h0e7: data <= 4'h6;
			10'h0e8: data <= 4'h7;
			10'h0e9: data <= 4'h1;
			10'h0ea: data <= 4'h0;
			10'h0eb: data <= 4'h4;
			10'h0ec: data <= 4'h2;
			10'h0ed: data <= 4'hd;
			10'h0ee: data <= 4'h0;
			10'h0ef: data <= 4'h0;
			10'h0f0: data <= 4'h1;
			10'h0f1: data <= 4'h8;
			10'h0f2: data <= 4'h0;
			10'h0f3: data <= 4'h0;
			10'h0f4: data <= 4'h8;
			10'h0f5: data <= 4'hc;
			10'h0f6: data <= 4'h3;
			10'h0f7: data <= 4'hb;
			10'h0f8: data <= 4'hd;
			10'h0f9: data <= 4'h3;
			10'h0fa: data <= 4'ha;
			10'h0fb: data <= 4'h1;
			10'h0fc: data <= 4'h3;
			10'h0fd: data <= 4'h5;
			10'h0fe: data <= 4'h6;
			10'h0ff: data <= 4'h5;
			10'h100: data <= 4'h6;
			10'h101: data <= 4'h5;
			10'h102: data <= 4'h6;
			10'h103: data <= 4'h5;
			10'h104: data <= 4'h5;
			10'h105: data <= 4'h6;
			10'h106: data <= 4'h6;
			10'h107: data <= 4'h5;
			10'h108: data <= 4'h6;
			10'h109: data <= 4'h6;
			10'h10a: data <= 4'h5;
			10'h10b: data <= 4'h5;
			10'h10c: data <= 4'h5;
			10'h10d: data <= 4'h4;
			10'h10e: data <= 4'h4;
			10'h10f: data <= 4'h6;
			10'h110: data <= 4'h6;
			10'h111: data <= 4'h7;
			10'h112: data <= 4'he;
			10'h113: data <= 4'h5;
			10'h114: data <= 4'h6;
			10'h115: data <= 4'h5;
			10'h116: data <= 4'h6;
			10'h117: data <= 4'h5;
			10'h118: data <= 4'h6;
			10'h119: data <= 4'h5;
			10'h11a: data <= 4'h5;
			10'h11b: data <= 4'h5;
			10'h11c: data <= 4'h6;
			10'h11d: data <= 4'h6;
			10'h11e: data <= 4'h6;
			10'h11f: data <= 4'h5;
			10'h120: data <= 4'h5;
			10'h121: data <= 4'h6;
			10'h122: data <= 4'h5;
			10'h123: data <= 4'h5;
			10'h124: data <= 4'h6;
			10'h125: data <= 4'h5;
			10'h126: data <= 4'h6;
			10'h127: data <= 4'h5;
			10'h128: data <= 4'h6;
			10'h129: data <= 4'h5;
			10'h12a: data <= 4'h6;
			10'h12b: data <= 4'h5;
			10'h12c: data <= 4'h6;
			10'h12d: data <= 4'h5;
			10'h12e: data <= 4'h5;
			10'h12f: data <= 4'h6;
			10'h130: data <= 4'h6;
			10'h131: data <= 4'h6;
			10'h132: data <= 4'h6;
			10'h133: data <= 4'h4;
			10'h134: data <= 4'h4;
			10'h135: data <= 4'h6;
			10'h136: data <= 4'h6;
			10'h137: data <= 4'h5;
			10'h138: data <= 4'h6;
			10'h139: data <= 4'h5;
			10'h13a: data <= 4'h6;
			10'h13b: data <= 4'h5;
			10'h13c: data <= 4'h6;
			10'h13d: data <= 4'h5;
			10'h13e: data <= 4'h5;
			10'h13f: data <= 4'h5;
			10'h140: data <= 4'h5;
			10'h141: data <= 4'h6;
			10'h142: data <= 4'h5;
			10'h143: data <= 4'h6;
			10'h144: data <= 4'h5;
			10'h145: data <= 4'h5;
			10'h146: data <= 4'h5;
			10'h147: data <= 4'h6;
			10'h148: data <= 4'h5;
			10'h149: data <= 4'h6;
			10'h14a: data <= 4'h5;
			10'h14b: data <= 4'h6;
			10'h14c: data <= 4'h5;
			10'h14d: data <= 4'h6;
			10'h14e: data <= 4'h5;
			10'h14f: data <= 4'h5;
			10'h150: data <= 4'h6;
			10'h151: data <= 4'h5;
			10'h152: data <= 4'h5;
			10'h153: data <= 4'h6;
			10'h154: data <= 4'h5;
			10'h155: data <= 4'h6;
			10'h156: data <= 4'h5;
			10'h157: data <= 4'h5;
			10'h158: data <= 4'h6;
			10'h159: data <= 4'h5;
			10'h15a: data <= 4'h6;
			10'h15b: data <= 4'h5;
			10'h15c: data <= 4'h6;
			10'h15d: data <= 4'h5;
			10'h15e: data <= 4'h6;
			10'h15f: data <= 4'h5;
			10'h160: data <= 4'h6;
			10'h161: data <= 4'h5;
			10'h162: data <= 4'h6;
			10'h163: data <= 4'h5;
			10'h164: data <= 4'h6;
			10'h165: data <= 4'h5;
			10'h166: data <= 4'h6;
			10'h167: data <= 4'h5;
			10'h168: data <= 4'h6;
			10'h169: data <= 4'h5;
			10'h16a: data <= 4'h6;
			10'h16b: data <= 4'h5;
			10'h16c: data <= 4'h6;
			10'h16d: data <= 4'h5;
			10'h16e: data <= 4'h6;
			10'h16f: data <= 4'h5;
			10'h170: data <= 4'h6;
			10'h171: data <= 4'h5;
			10'h172: data <= 4'h6;
			10'h173: data <= 4'h5;
			10'h174: data <= 4'h6;
			10'h175: data <= 4'h5;
			10'h176: data <= 4'h6;
			10'h177: data <= 4'h5;
			10'h178: data <= 4'h6;
			10'h179: data <= 4'h5;
			10'h17a: data <= 4'h6;
			10'h17b: data <= 4'h5;
			10'h17c: data <= 4'h6;
			10'h17d: data <= 4'h5;
			10'h17e: data <= 4'h6;
			10'h17f: data <= 4'h5;
			10'h180: data <= 4'h6;
			10'h181: data <= 4'h5;
			10'h182: data <= 4'h6;
			10'h183: data <= 4'h5;
			10'h184: data <= 4'h6;
			10'h185: data <= 4'h5;
			10'h186: data <= 4'h6;
			10'h187: data <= 4'h6;
			10'h188: data <= 4'h6;
			10'h189: data <= 4'h6;
			10'h18a: data <= 4'h5;
			10'h18b: data <= 4'h6;
			10'h18c: data <= 4'h6;
			10'h18d: data <= 4'h5;
			10'h18e: data <= 4'h6;
			10'h18f: data <= 4'h6;
			10'h190: data <= 4'h5;
			10'h191: data <= 4'h5;
			10'h192: data <= 4'h6;
			10'h193: data <= 4'h5;
			10'h194: data <= 4'h5;
			10'h195: data <= 4'h6;
			10'h196: data <= 4'h5;
			10'h197: data <= 4'h4;
			10'h198: data <= 4'h4;
			10'h199: data <= 4'h6;
			10'h19a: data <= 4'h6;
			10'h19b: data <= 4'h7;
			10'h19c: data <= 4'h1;
			10'h19d: data <= 4'h0;
			10'h19e: data <= 4'h4;
			10'h19f: data <= 4'h2;
			10'h1a0: data <= 4'hd;
			10'h1a1: data <= 4'h0;
			10'h1a2: data <= 4'h0;
			10'h1a3: data <= 4'h0;
			10'h1a4: data <= 4'h1;
			10'h1a5: data <= 4'h8;
			10'h1a6: data <= 4'h0;
			10'h1a7: data <= 4'h0;
			10'h1a8: data <= 4'h8;
			10'h1a9: data <= 4'h9;
			10'h1aa: data <= 4'h6;
			10'h1ab: data <= 4'hb;
			10'h1ac: data <= 4'ha;
			10'h1ad: data <= 4'h6;
			10'h1ae: data <= 4'h0;
			10'h1af: data <= 4'h0;
			10'h1b0: data <= 4'h5;
			10'h1b1: data <= 4'h6;
			10'h1b2: data <= 4'h5;
			10'h1b3: data <= 4'h6;
			10'h1b4: data <= 4'h5;
			10'h1b5: data <= 4'h6;
			10'h1b6: data <= 4'h5;
			10'h1b7: data <= 4'h5;
			10'h1b8: data <= 4'h5;
			10'h1b9: data <= 4'h6;
			10'h1ba: data <= 4'h5;
			10'h1bb: data <= 4'h5;
			10'h1bc: data <= 4'h6;
			10'h1bd: data <= 4'h6;
			10'h1be: data <= 4'h6;
			10'h1bf: data <= 4'h5;
			10'h1c0: data <= 4'h5;
			10'h1c1: data <= 4'h6;
			10'h1c2: data <= 4'h5;
			10'h1c3: data <= 4'h6;
			10'h1c4: data <= 4'h5;
			10'h1c5: data <= 4'h6;
			10'h1c6: data <= 4'h5;
			10'h1c7: data <= 4'h6;
			10'h1c8: data <= 4'h5;
			10'h1c9: data <= 4'h6;
			10'h1ca: data <= 4'h5;
			10'h1cb: data <= 4'h5;
			10'h1cc: data <= 4'h6;
			10'h1cd: data <= 4'h6;
			10'h1ce: data <= 4'h6;
			10'h1cf: data <= 4'h6;
			10'h1d0: data <= 4'h4;
			10'h1d1: data <= 4'h4;
			10'h1d2: data <= 4'h6;
			10'h1d3: data <= 4'h6;
			10'h1d4: data <= 4'h7;
			10'h1d5: data <= 4'h1;
			10'h1d6: data <= 4'h0;
			10'h1d7: data <= 4'h4;
			10'h1d8: data <= 4'h2;
			10'h1d9: data <= 4'hd;
			10'h1da: data <= 4'h0;
			10'h1db: data <= 4'h0;
			10'h1dc: data <= 4'h1;
			10'h1dd: data <= 4'h8;
			10'h1de: data <= 4'h0;
			10'h1df: data <= 4'h0;
			10'h1e0: data <= 4'h8;
			10'h1e1: data <= 4'h7;
			10'h1e2: data <= 4'h7;
			10'h1e3: data <= 4'hb;
			10'h1e4: data <= 4'h8;
			10'h1e5: data <= 4'h7;
			10'h1e6: data <= 4'ha;
			10'h1e7: data <= 4'hc;
			10'h1e8: data <= 4'h6;
			10'h1e9: data <= 4'h5;
			10'h1ea: data <= 4'h6;
			10'h1eb: data <= 4'h5;
			10'h1ec: data <= 4'h6;
			10'h1ed: data <= 4'h5;
			10'h1ee: data <= 4'h6;
			10'h1ef: data <= 4'h5;
			10'h1f0: data <= 4'h5;
			10'h1f1: data <= 4'h6;
			10'h1f2: data <= 4'h6;
			10'h1f3: data <= 4'h5;
			10'h1f4: data <= 4'h6;
			10'h1f5: data <= 4'h6;
			10'h1f6: data <= 4'h5;
			10'h1f7: data <= 4'h5;
			10'h1f8: data <= 4'h5;
			10'h1f9: data <= 4'h4;
			10'h1fa: data <= 4'h4;
			10'h1fb: data <= 4'h6;
			10'h1fc: data <= 4'h6;
			10'h1fd: data <= 4'h7;
			10'h1fe: data <= 4'hc;
			10'h1ff: data <= 4'h1;
			10'h200: data <= 4'h0;
			10'h201: data <= 4'h0;
			10'h202: data <= 4'hb;
			10'h203: data <= 4'h0;
			10'h204: data <= 4'h0;
			10'h205: data <= 4'h0;
			10'h206: data <= 4'h0;
			10'h207: data <= 4'h0;
			10'h208: data <= 4'h8;
			10'h209: data <= 4'ha;
			10'h20a: data <= 4'h9;
			10'h20b: data <= 4'h4;
			10'h20c: data <= 4'h4;
			10'h20d: data <= 4'h6;
			10'h20e: data <= 4'h6;
			10'h20f: data <= 4'h7;
			10'h210: data <= 4'hb;
			10'h211: data <= 4'h1;
			10'h212: data <= 4'h0;
			10'h213: data <= 4'he;
			10'h214: data <= 4'h5;
			10'h215: data <= 4'h6;
			10'h216: data <= 4'h5;
			10'h217: data <= 4'h6;
			10'h218: data <= 4'h5;
			10'h219: data <= 4'h6;
			10'h21a: data <= 4'h5;
			10'h21b: data <= 4'h5;
			10'h21c: data <= 4'h5;
			10'h21d: data <= 4'h6;
			10'h21e: data <= 4'h5;
			10'h21f: data <= 4'h5;
			10'h220: data <= 4'h6;
			10'h221: data <= 4'h6;
			10'h222: data <= 4'h6;
			10'h223: data <= 4'h5;
			10'h224: data <= 4'h5;
			10'h225: data <= 4'h6;
			10'h226: data <= 4'h5;
			10'h227: data <= 4'h6;
			10'h228: data <= 4'h5;
			10'h229: data <= 4'h6;
			10'h22a: data <= 4'h5;
			10'h22b: data <= 4'h5;
			10'h22c: data <= 4'h6;
			10'h22d: data <= 4'h5;
			10'h22e: data <= 4'h6;
			10'h22f: data <= 4'h6;
			10'h230: data <= 4'h6;
			10'h231: data <= 4'h5;
			10'h232: data <= 4'h5;
			10'h233: data <= 4'h6;
			10'h234: data <= 4'h4;
			10'h235: data <= 4'h4;
			10'h236: data <= 4'h6;
			10'h237: data <= 4'h6;
			10'h238: data <= 4'h7;
			10'h239: data <= 4'h1;
			10'h23a: data <= 4'h0;
			10'h23b: data <= 4'h4;
			10'h23c: data <= 4'h2;
			10'h23d: data <= 4'hd;
			10'h23e: data <= 4'h0;
			10'h23f: data <= 4'h0;
			10'h240: data <= 4'h1;
			10'h241: data <= 4'h8;
			10'h242: data <= 4'h0;
			10'h243: data <= 4'h0;
			10'h244: data <= 4'h8;
			10'h245: data <= 4'h0;
			10'h246: data <= 4'h9;
			10'h247: data <= 4'hb;
			10'h248: data <= 4'h1;
			10'h249: data <= 4'h9;
			10'h24a: data <= 4'ha;
			10'h24b: data <= 4'h0;
			10'h24c: data <= 4'h0;
			10'h24d: data <= 4'h5;
			10'h24e: data <= 4'h6;
			10'h24f: data <= 4'h5;
			10'h250: data <= 4'h6;
			10'h251: data <= 4'h5;
			10'h252: data <= 4'h6;
			10'h253: data <= 4'h5;
			10'h254: data <= 4'h5;
			10'h255: data <= 4'h6;
			10'h256: data <= 4'h6;
			10'h257: data <= 4'h5;
			10'h258: data <= 4'h6;
			10'h259: data <= 4'h6;
			10'h25a: data <= 4'h5;
			10'h25b: data <= 4'h5;
			10'h25c: data <= 4'h5;
			10'h25d: data <= 4'h4;
			10'h25e: data <= 4'h4;
			10'h25f: data <= 4'h6;
			10'h260: data <= 4'h6;
			10'h261: data <= 4'h7;
			10'h262: data <= 4'h1;
			10'h263: data <= 4'h0;
			10'h264: data <= 4'h0;
			10'h265: data <= 4'hb;
			10'h266: data <= 4'h0;
			10'h267: data <= 4'h0;
			10'h268: data <= 4'hc;
			10'h269: data <= 4'h1;
			10'h26a: data <= 4'h0;
			10'h26b: data <= 4'h0;
			10'h26c: data <= 4'hb;
			10'h26d: data <= 4'h0;
			10'h26e: data <= 4'h0;
			default: data <= 4'hX;
		endcase
	end
endmodule
